my name is humaira
my name is rehan 


