Hello!
Feature 1 added
