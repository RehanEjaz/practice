my name is humaira
